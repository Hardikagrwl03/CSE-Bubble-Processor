module instruction_memory(clk, rst, address, mode, write_data, out);

    input clk;
    input rst;
    input [4:0] address;
    input [31:0] write_data;
    input mode;
    output [31:0] out;

    reg [31:0] mem[24:0];
    reg [4:0] add_reg;
    reg [31:0] out;
    integer i = 1;

    initial begin
    mem[0] = 32'b00000000001000100000000000100000;
    mem[1] = 32'b00000000010000010000000000100010;
    mem[2] = 32'b00000000001000100000000000100001;
    mem[3] = 32'b00000000010000010000000000100011;
    mem[4] = 32'b00100000001000000000001111101000;
    mem[5] = 32'b00100100001000000000001111101000;
    mem[6] = 32'b00000000001000100000000000100100;
    mem[7] = 32'b00000000001000100000000000100101;
    mem[8] = 32'b00110000001000000000001111101000;
    mem[9] = 32'b00110100001000000000001111101000;
    mem[10] = 32'b00000000000000010000001010000000;
    mem[11] = 32'b00000000000000010000001010000010;
    mem[12] = 32'b10001100001000000000000000001010;
    mem[13] = 32'b10101100001000000000000000001010;
    mem[14] = 32'b00010000000000010000000000001010;
    mem[15] = 32'b00010100000000010000000000001010;
    mem[16] = 32'b00011100001000100000000000001010;
    mem[17] = 32'b00111100001000100000000000001010;
    mem[18] = 32'b00011000001000100000000000001010;
    mem[19] = 32'b01111100001000100000000000001010;
    mem[20] = 32'b00001000000000000000000000000010;
    mem[21] = 32'b00000000000000000000000000001000;
    mem[22] = 32'b00001100000000000000000000001010;
    mem[23] = 32'b00000000001000100000000000101010;
    mem[24] = 32'b00101000010000010000000001100100;
        
    end
    
    always @(posedge clk) begin
        add_reg <= address;
    end

    always @(mem[add_reg]) begin
        out <= mem[add_reg];
    end

    always @(posedge clk) begin
        if(mode == 1'b0)begin
            mem[address]=write_data;
        end
    end

    always @(posedge rst) begin
        mem[address] = 1'b0;
    end

endmodule